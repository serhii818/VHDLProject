

entity Uklad is
end Uklad;



architecture Uklad of Uklad is
begin



end Uklad;
