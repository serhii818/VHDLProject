
entity Uklad_tb is
end Uklad_tb;



architecture Uklad_tb of Uklad_tb is
begin



end Uklad_tb;
